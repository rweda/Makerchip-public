`line 2 "slide_example.m4out.tlv" 0

/*
Copyright (c) 2014, Intel Corporation

Redistribution and use in source and binary forms, with or without
modification, are permitted provided that the following conditions are met:

    * Redistributions of source code must retain the above copyright notice,
      this list of conditions and the following disclaimer.
    * Redistributions in binary form must reproduce the above copyright
      notice, this list of conditions and the following disclaimer in the
      documentation and/or other materials provided with the distribution.
    * Neither the name of Intel Corporation nor the names of its contributors
      may be used to endorse or promote products derived from this software
      without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE
FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/
   ...
// ---------- Generated Code Inlined Here (before 1st \TLV) ----------
`line 0 "slide_example.sv" 1
// Generated by SandPiper(TM).
// Redwood EDA, LLC does not claim intellectual property rights to this file and provides no warranty regarding its correctness or quality.


// For silencing unused signal messages.
`define BOGUS_USE(ignore)


genvar inst;


// Clock signals.
logic clkPV_sv_val ;

//
// Scope: |fetch
//

// For |fetch$valid.
logic FETCH_valid_a0;
logic FETCH_valid_a1;
logic FETCH_valid_a2;
logic FETCH_valid_a3;
logic FETCH_valid_a4;
logic FETCH_valid_a5;
logic FETCH_valid_a6;
logic FETCH_valid_a7;

// Clock signals.
logic clkP_FETCH_valid_a2 ;

//
// Scope: |fetch>inst[3:0]
//

// For |fetch>inst$g1_mem_op.
logic FETCH_Inst_g1_mem_op_a2 [3:0];
logic FETCH_Inst_g1_mem_op_a3 [3:0];
logic FETCH_Inst_g1_mem_op_a4 [3:0];
logic FETCH_Inst_g1_mem_op_a5 [3:0];
logic FETCH_Inst_g1_mem_op_a6 [3:0];

// For |fetch>inst$g3_immediate_op.
logic FETCH_Inst_g3_immediate_op_a2 [3:0];
logic FETCH_Inst_g3_immediate_op_a3 [3:0];
logic FETCH_Inst_g3_immediate_op_a4 [3:0];
logic FETCH_Inst_g3_immediate_op_a5 [3:0];
logic FETCH_Inst_g3_immediate_op_a6 [3:0];

// For |fetch>inst$immediate_op.
logic w_FETCH_Inst_immediate_op_a1 [3:0];
logic FETCH_Inst_immediate_op_a2 [3:0];

// For |fetch>inst$mem_op.
logic w_FETCH_Inst_mem_op_a1 [3:0];
logic FETCH_Inst_mem_op_a2 [3:0];

// For |fetch>inst$stuff1.
logic w_FETCH_Inst_stuff1_a2 [3:0];
logic FETCH_Inst_stuff1_a3 [3:0];
logic FETCH_Inst_stuff1_a4 [3:0];
logic FETCH_Inst_stuff1_a5 [3:0];
logic FETCH_Inst_stuff1_a6 [3:0];
logic FETCH_Inst_stuff1_a7 [3:0];

// For |fetch>inst$stuff2.
logic w_FETCH_Inst_stuff2_a2 [3:0];
logic FETCH_Inst_stuff2_a3 [3:0];
logic FETCH_Inst_stuff2_a4 [3:0];
logic FETCH_Inst_stuff2_a5 [3:0];
logic FETCH_Inst_stuff2_a6 [3:0];
logic FETCH_Inst_stuff2_a7 [3:0];

// Clock signals.
logic clkP_FETCH_Inst_g1_mem_op_a3 [3:0];
logic clkP_FETCH_Inst_g1_mem_op_a4 [3:0];
logic clkP_FETCH_Inst_g1_mem_op_a5 [3:0];
logic clkP_FETCH_Inst_g1_mem_op_a6 [3:0];
logic clkP_FETCH_Inst_g1_mem_op_a7 [3:0];
logic clkP_FETCH_Inst_g3_immediate_op_a3 [3:0];
logic clkP_FETCH_Inst_g3_immediate_op_a4 [3:0];
logic clkP_FETCH_Inst_g3_immediate_op_a5 [3:0];
logic clkP_FETCH_Inst_g3_immediate_op_a6 [3:0];
logic clkP_FETCH_Inst_g3_immediate_op_a7 [3:0];

//
// Scope: |pipe3
//

// For |pipe3$add.
logic PIPE3_add_a0;
logic PIPE3_add_a1;
logic PIPE3_add_a2;

// For |pipe3$best.
logic PIPE3_best_a1;
logic PIPE3_best_a2;
logic PIPE3_best_a3;
logic PIPE3_best_a4;
logic PIPE3_best_a5;

// For |pipe3$call.
logic PIPE3_call_a2;
logic PIPE3_call_a3;
logic PIPE3_call_a4;
logic PIPE3_call_a5;

// For |pipe3$git.
logic PIPE3_git_a5;
logic PIPE3_git_a6;
logic PIPE3_git_a7;
logic PIPE3_git_a8;
logic PIPE3_git_a9;
logic PIPE3_git_a10;
logic PIPE3_git_a11;

//
// Scope: |pipe6
//

//
// Scope: |pipe6>inst[3:0]
//

// For |pipe6>inst$mem_addr.
logic [50:0] w_PIPE6_Inst_mem_addr_a3L [3:0];
logic [50:0] PIPE6_Inst_mem_addr_a4L [3:0];

// For |pipe6>inst$mem_addr_plus1.
logic [50:0] PIPE6_Inst_mem_addr_plus1_a4L [3:0];

// For |pipe6>inst$raw_inst.
logic PIPE6_Inst_raw_inst_a1 [3:0];
logic PIPE6_Inst_raw_inst_a2 [3:0];
logic PIPE6_Inst_raw_inst_a3 [3:0];
logic PIPE6_Inst_raw_inst_a3L [3:0];

// For |pipe6>inst$valid.
logic PIPE6_Inst_valid_a0 [3:0];
logic PIPE6_Inst_valid_a1 [3:0];
logic PIPE6_Inst_valid_a2 [3:0];
logic PIPE6_Inst_valid_a3 [3:0];
logic PIPE6_Inst_valid_a3L [3:0];
logic PIPE6_Inst_valid_a4L [3:0];

// For |pipe6>inst$valid_mem_op.
logic w_PIPE6_Inst_valid_mem_op_a1 [3:0];

// Clock signals.
logic clkP_PIPE6_Inst_valid_a4L [3:0];

//
// Scope: |pipe7
//

// For |pipe7$foo.
logic PIPE7_foo_a1;



   //
   // Scope: |fetch
   //

      // Staging of $valid.
      always_ff @(posedge clk) FETCH_valid_a1 <= FETCH_valid_a0;
      always_ff @(posedge clk) FETCH_valid_a2 <= FETCH_valid_a1;
      always_ff @(posedge clk) FETCH_valid_a3 <= FETCH_valid_a2;
      always_ff @(posedge clk) FETCH_valid_a4 <= FETCH_valid_a3;
      always_ff @(posedge clk) FETCH_valid_a5 <= FETCH_valid_a4;
      always_ff @(posedge clk) FETCH_valid_a6 <= FETCH_valid_a5;
      always_ff @(posedge clk) FETCH_valid_a7 <= FETCH_valid_a6;


      //
      // Scope: >inst[3:0]
      //
      for (inst = 0; inst <= 3; inst++) begin : L1gen_FETCH_Inst
         // Staging of an unconditioned version of a condition signal.
         assign FETCH_Inst_g1_mem_op_a2[inst] = FETCH_Inst_mem_op_a2[inst] && FETCH_valid_a2;
         always_ff @(posedge clk) FETCH_Inst_g1_mem_op_a3[inst] <= FETCH_Inst_g1_mem_op_a2[inst];
         always_ff @(posedge clk) FETCH_Inst_g1_mem_op_a4[inst] <= FETCH_Inst_g1_mem_op_a3[inst];
         always_ff @(posedge clk) FETCH_Inst_g1_mem_op_a5[inst] <= FETCH_Inst_g1_mem_op_a4[inst];
         always_ff @(posedge clk) FETCH_Inst_g1_mem_op_a6[inst] <= FETCH_Inst_g1_mem_op_a5[inst];

         // Staging of an unconditioned version of a condition signal.
         assign FETCH_Inst_g3_immediate_op_a2[inst] = FETCH_Inst_immediate_op_a2[inst] && FETCH_valid_a2;
         always_ff @(posedge clk) FETCH_Inst_g3_immediate_op_a3[inst] <= FETCH_Inst_g3_immediate_op_a2[inst];
         always_ff @(posedge clk) FETCH_Inst_g3_immediate_op_a4[inst] <= FETCH_Inst_g3_immediate_op_a3[inst];
         always_ff @(posedge clk) FETCH_Inst_g3_immediate_op_a5[inst] <= FETCH_Inst_g3_immediate_op_a4[inst];
         always_ff @(posedge clk) FETCH_Inst_g3_immediate_op_a6[inst] <= FETCH_Inst_g3_immediate_op_a5[inst];

         // Staging of $immediate_op.
         always_ff @(posedge clkP_FETCH_valid_a2) FETCH_Inst_immediate_op_a2[inst] <= w_FETCH_Inst_immediate_op_a1[inst];

         // Staging of $mem_op.
         always_ff @(posedge clkP_FETCH_valid_a2) FETCH_Inst_mem_op_a2[inst] <= w_FETCH_Inst_mem_op_a1[inst];

         // Staging of $stuff1.
         always_ff @(posedge clkP_FETCH_Inst_g3_immediate_op_a3[inst]) FETCH_Inst_stuff1_a3[inst] <= w_FETCH_Inst_stuff1_a2[inst];
         always_ff @(posedge clkP_FETCH_Inst_g3_immediate_op_a4[inst]) FETCH_Inst_stuff1_a4[inst] <= FETCH_Inst_stuff1_a3[inst];
         always_ff @(posedge clkP_FETCH_Inst_g3_immediate_op_a5[inst]) FETCH_Inst_stuff1_a5[inst] <= FETCH_Inst_stuff1_a4[inst];
         always_ff @(posedge clkP_FETCH_Inst_g3_immediate_op_a6[inst]) FETCH_Inst_stuff1_a6[inst] <= FETCH_Inst_stuff1_a5[inst];
         always_ff @(posedge clkP_FETCH_Inst_g3_immediate_op_a7[inst]) FETCH_Inst_stuff1_a7[inst] <= FETCH_Inst_stuff1_a6[inst];

         // Staging of $stuff2.
         always_ff @(posedge clkP_FETCH_Inst_g1_mem_op_a3[inst]) FETCH_Inst_stuff2_a3[inst] <= w_FETCH_Inst_stuff2_a2[inst];
         always_ff @(posedge clkP_FETCH_Inst_g1_mem_op_a4[inst]) FETCH_Inst_stuff2_a4[inst] <= FETCH_Inst_stuff2_a3[inst];
         always_ff @(posedge clkP_FETCH_Inst_g1_mem_op_a5[inst]) FETCH_Inst_stuff2_a5[inst] <= FETCH_Inst_stuff2_a4[inst];
         always_ff @(posedge clkP_FETCH_Inst_g1_mem_op_a6[inst]) FETCH_Inst_stuff2_a6[inst] <= FETCH_Inst_stuff2_a5[inst];
         always_ff @(posedge clkP_FETCH_Inst_g1_mem_op_a7[inst]) FETCH_Inst_stuff2_a7[inst] <= FETCH_Inst_stuff2_a6[inst];

      end


   //
   // Scope: |pipe3
   //

      // Staging of $add.
      always_ff @(posedge clk) PIPE3_add_a1 <= PIPE3_add_a0;
      always_ff @(posedge clk) PIPE3_add_a2 <= PIPE3_add_a1;

      // Staging of $best.
      always_ff @(posedge clk) PIPE3_best_a2 <= PIPE3_best_a1;
      always_ff @(posedge clk) PIPE3_best_a3 <= PIPE3_best_a2;
      always_ff @(posedge clk) PIPE3_best_a4 <= PIPE3_best_a3;
      always_ff @(posedge clk) PIPE3_best_a5 <= PIPE3_best_a4;

      // Staging of $call.
      always_ff @(posedge clk) PIPE3_call_a3 <= PIPE3_call_a2;
      always_ff @(posedge clk) PIPE3_call_a4 <= PIPE3_call_a3;
      always_ff @(posedge clk) PIPE3_call_a5 <= PIPE3_call_a4;

      // Staging of $git.
      always_ff @(posedge clk) PIPE3_git_a6 <= PIPE3_git_a5;
      always_ff @(posedge clk) PIPE3_git_a7 <= PIPE3_git_a6;
      always_ff @(posedge clk) PIPE3_git_a8 <= PIPE3_git_a7;
      always_ff @(posedge clk) PIPE3_git_a9 <= PIPE3_git_a8;
      always_ff @(posedge clk) PIPE3_git_a10 <= PIPE3_git_a9;
      always_ff @(posedge clk) PIPE3_git_a11 <= PIPE3_git_a10;



   //
   // Scope: |pipe6
   //


      //
      // Scope: >inst[3:0]
      //
      for (inst = 0; inst <= 3; inst++) begin : L1gen_PIPE6_Inst
         // Staging of $mem_addr.
         always_ff @(posedge clkP_PIPE6_Inst_valid_a4L[inst]) PIPE6_Inst_mem_addr_a4L[inst][50:0] <= w_PIPE6_Inst_mem_addr_a3L[inst][50:0];

         // Staging of $raw_inst.
         always_ff @(posedge clkPV_sv_val) PIPE6_Inst_raw_inst_a2[inst] <= PIPE6_Inst_raw_inst_a1[inst];
         always_ff @(posedge clkPV_sv_val) PIPE6_Inst_raw_inst_a3[inst] <= PIPE6_Inst_raw_inst_a2[inst];
         always_latch if(clkPV_sv_val) PIPE6_Inst_raw_inst_a3L[inst] <= PIPE6_Inst_raw_inst_a3[inst];

         // Staging of $valid.
         always_ff @(posedge clk) PIPE6_Inst_valid_a1[inst] <= PIPE6_Inst_valid_a0[inst];
         always_ff @(posedge clk) PIPE6_Inst_valid_a2[inst] <= PIPE6_Inst_valid_a1[inst];
         always_ff @(posedge clk) PIPE6_Inst_valid_a3[inst] <= PIPE6_Inst_valid_a2[inst];
         always_latch if(n_clk) PIPE6_Inst_valid_a3L[inst] <= PIPE6_Inst_valid_a3[inst];
         always_ff @(posedge n_clk) PIPE6_Inst_valid_a4L[inst] <= PIPE6_Inst_valid_a3L[inst];

      end




//
// Gated clocks.
//


   clk_gate gen_clkPV_sv_val(clkPV_sv_val, clk, 1'b1, sv_val, 1'b0);

   //
   // Scope: |fetch
   //

      clk_gate gen_clkP_FETCH_valid_a2(clkP_FETCH_valid_a2, clk, 1'b1, FETCH_valid_a1, 1'b0);

      //
      // Scope: >inst[3:0]
      //
      for (inst = 0; inst <= 3; inst++) begin : L1clk_FETCH_Inst
         clk_gate gen_clkP_FETCH_Inst_g1_mem_op_a3(clkP_FETCH_Inst_g1_mem_op_a3[inst], clk, 1'b1, FETCH_Inst_g1_mem_op_a2[inst], 1'b0);
         clk_gate gen_clkP_FETCH_Inst_g1_mem_op_a4(clkP_FETCH_Inst_g1_mem_op_a4[inst], clk, 1'b1, FETCH_Inst_g1_mem_op_a3[inst], 1'b0);
         clk_gate gen_clkP_FETCH_Inst_g1_mem_op_a5(clkP_FETCH_Inst_g1_mem_op_a5[inst], clk, 1'b1, FETCH_Inst_g1_mem_op_a4[inst], 1'b0);
         clk_gate gen_clkP_FETCH_Inst_g1_mem_op_a6(clkP_FETCH_Inst_g1_mem_op_a6[inst], clk, 1'b1, FETCH_Inst_g1_mem_op_a5[inst], 1'b0);
         clk_gate gen_clkP_FETCH_Inst_g1_mem_op_a7(clkP_FETCH_Inst_g1_mem_op_a7[inst], clk, 1'b1, FETCH_Inst_g1_mem_op_a6[inst], 1'b0);
         clk_gate gen_clkP_FETCH_Inst_g3_immediate_op_a3(clkP_FETCH_Inst_g3_immediate_op_a3[inst], clk, 1'b1, FETCH_Inst_g3_immediate_op_a2[inst], 1'b0);
         clk_gate gen_clkP_FETCH_Inst_g3_immediate_op_a4(clkP_FETCH_Inst_g3_immediate_op_a4[inst], clk, 1'b1, FETCH_Inst_g3_immediate_op_a3[inst], 1'b0);
         clk_gate gen_clkP_FETCH_Inst_g3_immediate_op_a5(clkP_FETCH_Inst_g3_immediate_op_a5[inst], clk, 1'b1, FETCH_Inst_g3_immediate_op_a4[inst], 1'b0);
         clk_gate gen_clkP_FETCH_Inst_g3_immediate_op_a6(clkP_FETCH_Inst_g3_immediate_op_a6[inst], clk, 1'b1, FETCH_Inst_g3_immediate_op_a5[inst], 1'b0);
         clk_gate gen_clkP_FETCH_Inst_g3_immediate_op_a7(clkP_FETCH_Inst_g3_immediate_op_a7[inst], clk, 1'b1, FETCH_Inst_g3_immediate_op_a6[inst], 1'b0);
      end


   //
   // Scope: |pipe6
   //


      //
      // Scope: >inst[3:0]
      //
      for (inst = 0; inst <= 3; inst++) begin : L1clk_PIPE6_Inst
         clk_gate gen_clkP_PIPE6_Inst_valid_a4L(clkP_PIPE6_Inst_valid_a4L[inst], n_clk, 1'b1, PIPE6_Inst_valid_a3L[inst], 1'b0);
      end


// ---------- Generated Code Ends ----------
`line 32 "slide_example.m4out.tlv"
//_\TLV
   //_|fetch
      //_@0
         assign FETCH_valid_a0 = stuff;
      //_?$valid
         for (inst = 0; inst <= 3; inst++) begin : L1_FETCH_Inst //_>inst
            //_@1
               assign w_FETCH_Inst_mem_op_a1[inst] = decode;
               assign w_FETCH_Inst_immediate_op_a1[inst] = decode;
            //_?$mem_op
               //_?$immediate_op
                  //_@2
                     assign w_FETCH_Inst_stuff1_a2[inst] = exp;
            //_?$immediate_op
               //_?$mem_op
                  //_@2
                     assign w_FETCH_Inst_stuff2_a2[inst] = exp;
            //_@7
               `BOGUS_USE(FETCH_Inst_stuff1_a7[inst], FETCH_Inst_stuff2_a7[inst]) end
   //_|pipe6
      //@0
      //   $blah = stuff3;
      for (inst = 0; inst <= 3; inst++) begin : L1_PIPE6_Inst //_>inst
         //_@0
            assign PIPE6_Inst_valid_a0[inst] = valid_U600H;
            assign sv_val = stuff4;
         //_?*sv_val
            //_@1
               assign PIPE6_Inst_raw_inst_a1[inst] = ...;
               assign w_PIPE6_Inst_valid_mem_op_a1[inst] = PIPE6_Inst_raw_inst_a1[inst] == 2'b01;
            //_?$valid
               //_@3.1
                  assign w_PIPE6_Inst_mem_addr_a3L[inst][50:0] = /*$op_a +*/ PIPE6_Inst_raw_inst_a3L[inst];
               //_@4.1
                  assign PIPE6_Inst_mem_addr_plus1_a4L[inst][50:0] = PIPE6_Inst_mem_addr_a4L[inst] | 51'b1;   // BUG: Enable for the clock producing $mem_addr@4L is not created.
                  `BOGUS_USE(PIPE6_Inst_mem_addr_plus1_a4L[inst]) end
   //_|pipe7
      //_@1
         assign PIPE7_foo_a1 = PIPE6_Inst_valid_a1[0];
         `BOGUS_USE(PIPE7_foo_a1)
   //_|pipe3
      //_@0
         assign PIPE3_add_a0 = valid_U400H;
      //_@1
         assign PIPE3_best_a1 = PIPE3_add_a1;
      //_@2
         assign PIPE3_call_a2 = PIPE3_add_a2 | PIPE3_best_a2;
      //_@5
         assign PIPE3_git_a5 = PIPE3_call_a5 | PIPE3_best_a5;
   //_|pipe4
      //_@1
         `MACRO(PIPE3_add_a0 + PIPE3_git_a11)



// Undefine macros defined by SandPiper.
`undef BOGUS_USE
