`line 2 "ring.m4out.tlv" 0

/*
Copyright (c) 2014, Intel Corporation

Redistribution and use in source and binary forms, with or without
modification, are permitted provided that the following conditions are met:

    * Redistributions of source code must retain the above copyright notice,
      this list of conditions and the following disclaimer.
    * Redistributions in binary form must reproduce the above copyright
      notice, this list of conditions and the following disclaimer in the
      documentation and/or other materials provided with the distribution.
    * Neither the name of Intel Corporation nor the names of its contributors
      may be used to endorse or promote products derived from this software
      without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE
FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

`include "ring.vh"



module ring (
   // Primary inputs
   input logic clk,
   input logic reset,

   input logic [7:0] data_in [RING_STOPS],
   input logic [RING_STOPS_WIDTH-1:0] dest_in [RING_STOPS],
   input logic valid_in [RING_STOPS],

   // Primary outputs
   output logic accepted [RING_STOPS],
   output logic [7:0] data_out [RING_STOPS],
   output logic valid_out [RING_STOPS]
);

// ---------- Generated Code Inlined Here (before 1st \TLV) ----------
`line 0 "ring.sv" 1
// Generated by SandPiper(TM).
// Redwood EDA, LLC does not claim intellectual property rights to this file and provides no warranty regarding its correctness or quality.


// For silencing unused signal messages.
`define BOGUS_USE(ignore)


// For X injection on assignments, disableable using `define SP_PHYS.
`ifdef WHEN
   $warning("WHEN macro redefined.");
`endif
`ifdef SP_PHYS
   `define WHEN(valid_sig)
`else
   `define WHEN(valid_sig) !valid_sig ? 'x :
`endif


genvar entry, stop;


//
// Scope: >stop[RING_STOPS-1:0]
//

//
// Scope: >stop|fo
//

// For >stop|fo$blocked.
logic [RING_STOPS-1:0] Stop_FO_blocked_a0;

// For >stop|fo$data.
logic [RING_STOPS-1:0] [7:0] w_Stop_FO_data_a0 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] [7:0] Stop_FO_data_a0;
logic [RING_STOPS-1:0] [7:0] Stop_FO_data_a1;

// For >stop|fo$dest.
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] w_Stop_FO_dest_a0 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] Stop_FO_dest_a0;

// For >stop|fo$parity.
logic [RING_STOPS-1:0] w_Stop_FO_parity_a0 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] Stop_FO_parity_a0;
logic [RING_STOPS-1:0] Stop_FO_parity_a1;

// For >stop|fo$trans_avail.
logic [RING_STOPS-1:0] Stop_FO_trans_avail_a0;

// For >stop|fo$trans_valid.
logic [RING_STOPS-1:0] Stop_FO_trans_valid_a0;

// Clock signals.
logic clkP_Stop_FO_trans_valid_a1 [RING_STOPS-1:0];

//
// Scope: >stop|fo>entry[(6)-1:0]
//

// For >stop|fo>entry$is_head.
logic [RING_STOPS-1:0][(6)-1:0] Stop_FO_Entry_is_head_a0;

// For >stop|fo>entry$pop.
logic [RING_STOPS-1:0][(6)-1:0] Stop_FO_Entry_pop_a0;

//
// Scope: >stop|fo>entry>accum
//

// For >stop|fo>entry>accum$data.
logic [RING_STOPS-1:0][(6)-1:0] [7:0] Stop_FO_Entry_Accum_data_a0;

// For >stop|fo>entry>accum$dest.
logic [RING_STOPS-1:0][(6)-1:0] [RING_STOPS_WIDTH-1:0] Stop_FO_Entry_Accum_dest_a0;

// For >stop|fo>entry>accum$parity.
logic [RING_STOPS-1:0][(6)-1:0] Stop_FO_Entry_Accum_parity_a0;

//
// Scope: >stop|fo>entry>read_masked
//

// For >stop|fo>entry>read_masked$data.
logic [RING_STOPS-1:0][(6)-1:0] [7:0] Stop_FO_Entry_ReadMasked_data_a0;

// For >stop|fo>entry>read_masked$dest.
logic [RING_STOPS-1:0][(6)-1:0] [RING_STOPS_WIDTH-1:0] Stop_FO_Entry_ReadMasked_dest_a0;

// For >stop|fo>entry>read_masked$parity.
logic [RING_STOPS-1:0][(6)-1:0] Stop_FO_Entry_ReadMasked_parity_a0;

//
// Scope: >stop|fo>fifo_head
//

// For >stop|fo>fifo_head$data.
logic [RING_STOPS-1:0] [7:0] w_Stop_FO_FifoHead_data_a0 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] [7:0] Stop_FO_FifoHead_data_a0;

// For >stop|fo>fifo_head$dest.
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] w_Stop_FO_FifoHead_dest_a0 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] Stop_FO_FifoHead_dest_a0;

// For >stop|fo>fifo_head$parity.
logic [RING_STOPS-1:0] w_Stop_FO_FifoHead_parity_a0 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] Stop_FO_FifoHead_parity_a0;

// For >stop|fo>fifo_head$trans_avail.
logic [RING_STOPS-1:0] Stop_FO_FifoHead_trans_avail_a0;

//
// Scope: >stop|fo>head
//

// For >stop|fo>head$data.
logic [RING_STOPS-1:0] [7:0] w_Stop_FO_Head_data_a0 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] [7:0] Stop_FO_Head_data_a0;

// For >stop|fo>head$dest.
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] w_Stop_FO_Head_dest_a0 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] Stop_FO_Head_dest_a0;

// For >stop|fo>head$parity.
logic [RING_STOPS-1:0] w_Stop_FO_Head_parity_a0 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] Stop_FO_Head_parity_a0;

// For >stop|fo>head$trans_avail.
logic [RING_STOPS-1:0] Stop_FO_Head_trans_avail_a0;

//
// Scope: >stop|inpipe
//

// For >stop|inpipe$blocked.
logic [RING_STOPS-1:0] Stop_INPIPE_blocked_a1;

// For >stop|inpipe$bypass.
logic [RING_STOPS-1:0] Stop_INPIPE_bypass_a1;

// For >stop|inpipe$data.
logic [RING_STOPS-1:0] [7:0] Stop_INPIPE_data_a0;
logic [RING_STOPS-1:0] [7:0] Stop_INPIPE_data_a1;

// For >stop|inpipe$dest.
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] Stop_INPIPE_dest_a0;
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] Stop_INPIPE_dest_a1;

// For >stop|inpipe$empty.
logic [RING_STOPS-1:0] Stop_INPIPE_empty_a2;

// For >stop|inpipe$full.
logic [RING_STOPS-1:0] Stop_INPIPE_full_a2;

// For >stop|inpipe$grow.
logic [RING_STOPS-1:0] Stop_INPIPE_grow_a1;

// For >stop|inpipe$out_blocked.
logic [RING_STOPS-1:0] Stop_INPIPE_out_blocked_a1;

// For >stop|inpipe$parity.
logic [RING_STOPS-1:0] Stop_INPIPE_parity_a0;
logic [RING_STOPS-1:0] Stop_INPIPE_parity_a1;

// For >stop|inpipe$push.
logic [RING_STOPS-1:0] Stop_INPIPE_push_a1;

// For >stop|inpipe$reset.
logic [RING_STOPS-1:0] Stop_INPIPE_reset_a1;

// For >stop|inpipe$shrink.
logic [RING_STOPS-1:0] Stop_INPIPE_shrink_a1;

// For >stop|inpipe$trans_avail.
logic [RING_STOPS-1:0] Stop_INPIPE_trans_avail_a0;
logic [RING_STOPS-1:0] Stop_INPIPE_trans_avail_a1;

// For >stop|inpipe$trans_valid.
logic [RING_STOPS-1:0] Stop_INPIPE_trans_valid_a1;

// For >stop|inpipe$two_valid.
logic [RING_STOPS-1:0] Stop_INPIPE_two_valid_a1;
logic [RING_STOPS-1:0] Stop_INPIPE_two_valid_a2;

// For >stop|inpipe$valid_count.
logic [RING_STOPS-1:0] [$clog2((6)+1)-1:0] Stop_INPIPE_valid_count_a1;
logic [RING_STOPS-1:0] [$clog2((6)+1)-1:0] Stop_INPIPE_valid_count_a2;

// For >stop|inpipe$would_bypass.
logic [RING_STOPS-1:0] Stop_INPIPE_would_bypass_a1;

//
// Scope: >stop|inpipe>entry[(6)-1:0]
//

// For >stop|inpipe>entry$State.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_State_a1;
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_State_a2;

// For >stop|inpipe>entry$data.
logic [RING_STOPS-1:0][(6)-1:0] [7:0] Stop_INPIPE_Entry_data_a1;
logic [RING_STOPS-1:0][(6)-1:0] [7:0] Stop_INPIPE_Entry_data_a2;

// For >stop|inpipe>entry$dest.
logic [RING_STOPS-1:0][(6)-1:0] [RING_STOPS_WIDTH-1:0] Stop_INPIPE_Entry_dest_a1;
logic [RING_STOPS-1:0][(6)-1:0] [RING_STOPS_WIDTH-1:0] Stop_INPIPE_Entry_dest_a2;

// For >stop|inpipe>entry$is_head.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_is_head_a2;

// For >stop|inpipe>entry$is_tail.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_is_tail_a1;

// For >stop|inpipe>entry$next_entry_state.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_next_entry_state_a2;

// For >stop|inpipe>entry$parity.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_parity_a1;
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_parity_a2;

// For >stop|inpipe>entry$prev_entry_state.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_prev_entry_state_a2;

// For >stop|inpipe>entry$prev_entry_was_tail.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_prev_entry_was_tail_a1;

// For >stop|inpipe>entry$push.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_push_a1;

// For >stop|inpipe>entry$reconstructed_is_tail.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_reconstructed_is_tail_a2;

// For >stop|inpipe>entry$reconstructed_valid.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_reconstructed_valid_a2;

// For >stop|inpipe>entry$valid.
logic [RING_STOPS-1:0][(6)-1:0] Stop_INPIPE_Entry_valid_a1;

//
// Scope: >stop|outpipe
//

// For >stop|outpipe$blocked.
logic [RING_STOPS-1:0] Stop_OUTPIPE_blocked_a0;

// For >stop|outpipe$data.
logic [RING_STOPS-1:0] [7:0] w_Stop_OUTPIPE_data_a1 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] [7:0] Stop_OUTPIPE_data_a1;
logic [RING_STOPS-1:0] [7:0] Stop_OUTPIPE_data_a2;

// For >stop|outpipe$parity.
logic [RING_STOPS-1:0] w_Stop_OUTPIPE_parity_a1 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] Stop_OUTPIPE_parity_a1;
logic [RING_STOPS-1:0] Stop_OUTPIPE_parity_a2;

// For >stop|outpipe$trans_avail.
logic [RING_STOPS-1:0] Stop_OUTPIPE_trans_avail_a0;

// For >stop|outpipe$trans_valid.
logic [RING_STOPS-1:0] Stop_OUTPIPE_trans_valid_a0;
logic [RING_STOPS-1:0] Stop_OUTPIPE_trans_valid_a1;
logic [RING_STOPS-1:0] Stop_OUTPIPE_trans_valid_a2;

// Clock signals.
logic clkP_Stop_OUTPIPE_trans_valid_a2 [RING_STOPS-1:0];

//
// Scope: >stop|rg
//

// For >stop|rg$data.
logic [RING_STOPS-1:0] [7:0] w_Stop_RG_data_a1 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] [7:0] Stop_RG_data_a1;
logic [RING_STOPS-1:0] [7:0] Stop_RG_data_a2;

// For >stop|rg$dest.
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] Stop_RG_dest_a0;
logic [RING_STOPS-1:0] [RING_STOPS_WIDTH-1:0] Stop_RG_dest_a1;

// For >stop|rg$parity.
logic [RING_STOPS-1:0] w_Stop_RG_parity_a1 /* without X injection for "when" condition */;
logic [RING_STOPS-1:0] Stop_RG_parity_a1;
logic [RING_STOPS-1:0] Stop_RG_parity_a2;

// For >stop|rg$pass_on.
logic [RING_STOPS-1:0] Stop_RG_pass_on_a0;
logic [RING_STOPS-1:0] Stop_RG_pass_on_a1;

// For >stop|rg$passed_on.
logic [RING_STOPS-1:0] Stop_RG_passed_on_a0;
logic [RING_STOPS-1:0] Stop_RG_passed_on_a1;

// For >stop|rg$valid.
logic [RING_STOPS-1:0] Stop_RG_valid_a0;
logic [RING_STOPS-1:0] Stop_RG_valid_a1;

// Clock signals.
logic clkP_Stop_RG_valid_a2 [RING_STOPS-1:0];

//
// Scope: |reset
//

// For |reset$reset.
logic RESET_reset_a0;
logic RESET_reset_a1;
logic RESET_reset_a2;



   //
   // Scope: >stop[RING_STOPS-1:0]
   //
   for (stop = 0; stop <= RING_STOPS-1; stop++) begin : L1gen_Stop

      //
      // Scope: |fo
      //

         // Inject X when invalid.
         assign Stop_FO_data_a0[stop] = `WHEN(Stop_FO_trans_valid_a0[stop]) w_Stop_FO_data_a0[stop];
         // Staging of $data.
         always_ff @(posedge clkP_Stop_FO_trans_valid_a1[stop]) Stop_FO_data_a1[stop][7:0] <= Stop_FO_data_a0[stop][7:0];

         // Inject X when invalid.
         assign Stop_FO_dest_a0[stop] = `WHEN(Stop_FO_trans_valid_a0[stop]) w_Stop_FO_dest_a0[stop];
         // Inject X when invalid.
         assign Stop_FO_parity_a0[stop] = `WHEN(Stop_FO_trans_valid_a0[stop]) w_Stop_FO_parity_a0[stop];
         // Staging of $parity.
         always_ff @(posedge clkP_Stop_FO_trans_valid_a1[stop]) Stop_FO_parity_a1[stop] <= Stop_FO_parity_a0[stop];


         //
         // Scope: >fifo_head
         //

            // Inject X when invalid.
            assign Stop_FO_FifoHead_data_a0[stop] = `WHEN(Stop_FO_FifoHead_trans_avail_a0[stop]) w_Stop_FO_FifoHead_data_a0[stop];
            // Inject X when invalid.
            assign Stop_FO_FifoHead_dest_a0[stop] = `WHEN(Stop_FO_FifoHead_trans_avail_a0[stop]) w_Stop_FO_FifoHead_dest_a0[stop];
            // Inject X when invalid.
            assign Stop_FO_FifoHead_parity_a0[stop] = `WHEN(Stop_FO_FifoHead_trans_avail_a0[stop]) w_Stop_FO_FifoHead_parity_a0[stop];


         //
         // Scope: >head
         //

            // Inject X when invalid.
            assign Stop_FO_Head_data_a0[stop] = `WHEN(Stop_FO_Head_trans_avail_a0[stop]) w_Stop_FO_Head_data_a0[stop];
            // Inject X when invalid.
            assign Stop_FO_Head_dest_a0[stop] = `WHEN(Stop_FO_Head_trans_avail_a0[stop]) w_Stop_FO_Head_dest_a0[stop];
            // Inject X when invalid.
            assign Stop_FO_Head_parity_a0[stop] = `WHEN(Stop_FO_Head_trans_avail_a0[stop]) w_Stop_FO_Head_parity_a0[stop];



      //
      // Scope: |inpipe
      //

         // Staging of $data.
         always_ff @(posedge clk) Stop_INPIPE_data_a1[stop][7:0] <= Stop_INPIPE_data_a0[stop][7:0];

         // Staging of $dest.
         always_ff @(posedge clk) Stop_INPIPE_dest_a1[stop][RING_STOPS_WIDTH-1:0] <= Stop_INPIPE_dest_a0[stop][RING_STOPS_WIDTH-1:0];

         // Staging of $parity.
         always_ff @(posedge clk) Stop_INPIPE_parity_a1[stop] <= Stop_INPIPE_parity_a0[stop];

         // Staging of $trans_avail.
         always_ff @(posedge clk) Stop_INPIPE_trans_avail_a1[stop] <= Stop_INPIPE_trans_avail_a0[stop];

         // Staging of $two_valid.
         always_ff @(posedge clk) Stop_INPIPE_two_valid_a2[stop] <= Stop_INPIPE_two_valid_a1[stop];

         // Staging of $valid_count.
         always_ff @(posedge clk) Stop_INPIPE_valid_count_a2[stop][$clog2((6)+1)-1:0] <= Stop_INPIPE_valid_count_a1[stop][$clog2((6)+1)-1:0];


         //
         // Scope: >entry[(6)-1:0]
         //
         for (entry = 0; entry <= (6)-1; entry++) begin : L2gen_INPIPE_Entry
            // Staging of $State.
            always_ff @(posedge clk) Stop_INPIPE_Entry_State_a2[stop][entry] <= Stop_INPIPE_Entry_State_a1[stop][entry];

            // Staging of $data.
            always_ff @(posedge clk) Stop_INPIPE_Entry_data_a2[stop][entry][7:0] <= Stop_INPIPE_Entry_data_a1[stop][entry][7:0];

            // Staging of $dest.
            always_ff @(posedge clk) Stop_INPIPE_Entry_dest_a2[stop][entry][RING_STOPS_WIDTH-1:0] <= Stop_INPIPE_Entry_dest_a1[stop][entry][RING_STOPS_WIDTH-1:0];

            // Staging of $parity.
            always_ff @(posedge clk) Stop_INPIPE_Entry_parity_a2[stop][entry] <= Stop_INPIPE_Entry_parity_a1[stop][entry];

         end


      //
      // Scope: |outpipe
      //

         // Inject X when invalid.
         assign Stop_OUTPIPE_data_a1[stop] = `WHEN(Stop_OUTPIPE_trans_valid_a1[stop]) w_Stop_OUTPIPE_data_a1[stop];
         // Staging of $data.
         always_ff @(posedge clkP_Stop_OUTPIPE_trans_valid_a2[stop]) Stop_OUTPIPE_data_a2[stop][7:0] <= Stop_OUTPIPE_data_a1[stop][7:0];

         // Inject X when invalid.
         assign Stop_OUTPIPE_parity_a1[stop] = `WHEN(Stop_OUTPIPE_trans_valid_a1[stop]) w_Stop_OUTPIPE_parity_a1[stop];
         // Staging of $parity.
         always_ff @(posedge clkP_Stop_OUTPIPE_trans_valid_a2[stop]) Stop_OUTPIPE_parity_a2[stop] <= Stop_OUTPIPE_parity_a1[stop];

         // Staging of $trans_valid.
         always_ff @(posedge clk) Stop_OUTPIPE_trans_valid_a1[stop] <= Stop_OUTPIPE_trans_valid_a0[stop];
         always_ff @(posedge clk) Stop_OUTPIPE_trans_valid_a2[stop] <= Stop_OUTPIPE_trans_valid_a1[stop];



      //
      // Scope: |rg
      //

         // Inject X when invalid.
         assign Stop_RG_data_a1[stop] = `WHEN(Stop_RG_valid_a1[stop]) w_Stop_RG_data_a1[stop];
         // Staging of $data.
         always_ff @(posedge clkP_Stop_RG_valid_a2[stop]) Stop_RG_data_a2[stop][7:0] <= Stop_RG_data_a1[stop][7:0];

         // Staging of $dest.
         always_ff @(posedge clk) Stop_RG_dest_a1[stop][RING_STOPS_WIDTH-1:0] <= Stop_RG_dest_a0[stop][RING_STOPS_WIDTH-1:0];

         // Inject X when invalid.
         assign Stop_RG_parity_a1[stop] = `WHEN(Stop_RG_valid_a1[stop]) w_Stop_RG_parity_a1[stop];
         // Staging of $parity.
         always_ff @(posedge clkP_Stop_RG_valid_a2[stop]) Stop_RG_parity_a2[stop] <= Stop_RG_parity_a1[stop];

         // Staging of $pass_on.
         always_ff @(posedge clk) Stop_RG_pass_on_a1[stop] <= Stop_RG_pass_on_a0[stop];

         // Staging of $passed_on.
         always_ff @(posedge clk) Stop_RG_passed_on_a1[stop] <= Stop_RG_passed_on_a0[stop];

         // Staging of $valid.
         always_ff @(posedge clk) Stop_RG_valid_a1[stop] <= Stop_RG_valid_a0[stop];


   end

   //
   // Scope: |reset
   //

      // Staging of $reset.
      always_ff @(posedge clk) RESET_reset_a1 <= RESET_reset_a0;
      always_ff @(posedge clk) RESET_reset_a2 <= RESET_reset_a1;





//
// Gated clocks.
//



   //
   // Scope: >stop[RING_STOPS-1:0]
   //
   for (stop = 0; stop <= RING_STOPS-1; stop++) begin : L1clk_Stop

      //
      // Scope: |fo
      //

         clk_gate gen_clkP_Stop_FO_trans_valid_a1(clkP_Stop_FO_trans_valid_a1[stop], clk, 1'b1, (Stop_FO_trans_valid_a0[stop] ? 1'b1 : 1'bx), 1'b0);


      //
      // Scope: |outpipe
      //

         clk_gate gen_clkP_Stop_OUTPIPE_trans_valid_a2(clkP_Stop_OUTPIPE_trans_valid_a2[stop], clk, 1'b1, (Stop_OUTPIPE_trans_valid_a1[stop] ? 1'b1 : 1'bx), 1'b0);


      //
      // Scope: |rg
      //

         clk_gate gen_clkP_Stop_RG_valid_a2(clkP_Stop_RG_valid_a2[stop], clk, 1'b1, (Stop_RG_valid_a1[stop] ? 1'b1 : 1'bx), 1'b0);

   end




//
// Debug Signals
//

   if (1) begin : DEBUG_SIGS


      //
      // Scope: >stop[RING_STOPS-1:0]
      //
      for (stop = 0; stop <= RING_STOPS-1; stop++) begin : \>stop 

         //
         // Scope: |fo
         //
         if (1) begin : \|fo 
            logic  \//?$trans_valid@0$ANY ;
            assign \//?$trans_valid@0$ANY  = 1'b1;
            logic  \//@0$blocked ;
            assign \//@0$blocked = Stop_FO_blocked_a0[stop];
            logic [7:0] \//?$trans_valid@0$data ;
            assign \//?$trans_valid@0$data = Stop_FO_data_a0[stop];
            logic [RING_STOPS_WIDTH-1:0] \//?$trans_valid@0$dest ;
            assign \//?$trans_valid@0$dest = Stop_FO_dest_a0[stop];
            logic  \//?$trans_valid@0$parity ;
            assign \//?$trans_valid@0$parity = Stop_FO_parity_a0[stop];
            logic  \//@0$trans_avail ;
            assign \//@0$trans_avail = Stop_FO_trans_avail_a0[stop];
            logic  \//@0$trans_valid ;
            assign \//@0$trans_valid = Stop_FO_trans_valid_a0[stop];

            //
            // Scope: >entry[(6)-1:0]
            //
            for (entry = 0; entry <= (6)-1; entry++) begin : \>entry 
               logic  \///@0$is_head ;
               assign \///@0$is_head = Stop_FO_Entry_is_head_a0[stop][entry];
               logic  \///@0$pop ;
               assign \///@0$pop = Stop_FO_Entry_pop_a0[stop][entry];

               //
               // Scope: >accum
               //
               if (1) begin : \>accum 
                  logic  \////@0$ANY ;
                  assign \////@0$ANY  = 1'b1;
                  logic [7:0] \////@0$data ;
                  assign \////@0$data = Stop_FO_Entry_Accum_data_a0[stop][entry];
                  logic [RING_STOPS_WIDTH-1:0] \////@0$dest ;
                  assign \////@0$dest = Stop_FO_Entry_Accum_dest_a0[stop][entry];
                  logic  \////@0$parity ;
                  assign \////@0$parity = Stop_FO_Entry_Accum_parity_a0[stop][entry];
               end

               //
               // Scope: >read_masked
               //
               if (1) begin : \>read_masked 
                  logic  \////@0$ANY ;
                  assign \////@0$ANY  = 1'b1;
                  logic [7:0] \////@0$data ;
                  assign \////@0$data = Stop_FO_Entry_ReadMasked_data_a0[stop][entry];
                  logic [RING_STOPS_WIDTH-1:0] \////@0$dest ;
                  assign \////@0$dest = Stop_FO_Entry_ReadMasked_dest_a0[stop][entry];
                  logic  \////@0$parity ;
                  assign \////@0$parity = Stop_FO_Entry_ReadMasked_parity_a0[stop][entry];
               end
            end

            //
            // Scope: >fifo_head
            //
            if (1) begin : \>fifo_head 
               logic  \///?$trans_avail@0$ANY ;
               assign \///?$trans_avail@0$ANY  = 1'b1;
               logic [7:0] \///?$trans_avail@0$data ;
               assign \///?$trans_avail@0$data = Stop_FO_FifoHead_data_a0[stop];
               logic [RING_STOPS_WIDTH-1:0] \///?$trans_avail@0$dest ;
               assign \///?$trans_avail@0$dest = Stop_FO_FifoHead_dest_a0[stop];
               logic  \///?$trans_avail@0$parity ;
               assign \///?$trans_avail@0$parity = Stop_FO_FifoHead_parity_a0[stop];
               logic  \///@0$trans_avail ;
               assign \///@0$trans_avail = Stop_FO_FifoHead_trans_avail_a0[stop];
            end

            //
            // Scope: >head
            //
            if (1) begin : \>head 
               logic  \///?$trans_avail@0$ANY ;
               assign \///?$trans_avail@0$ANY  = 1'b1;
               logic [7:0] \///?$trans_avail@0$data ;
               assign \///?$trans_avail@0$data = Stop_FO_Head_data_a0[stop];
               logic [RING_STOPS_WIDTH-1:0] \///?$trans_avail@0$dest ;
               assign \///?$trans_avail@0$dest = Stop_FO_Head_dest_a0[stop];
               logic  \///?$trans_avail@0$parity ;
               assign \///?$trans_avail@0$parity = Stop_FO_Head_parity_a0[stop];
               logic  \///@0$trans_avail ;
               assign \///@0$trans_avail = Stop_FO_Head_trans_avail_a0[stop];
            end
         end

         //
         // Scope: |inpipe
         //
         if (1) begin : \|inpipe 
            logic  \//@1$blocked ;
            assign \//@1$blocked = Stop_INPIPE_blocked_a1[stop];
            logic  \//@1$bypass ;
            assign \//@1$bypass = Stop_INPIPE_bypass_a1[stop];
            logic [7:0] \//@0$data ;
            assign \//@0$data = Stop_INPIPE_data_a0[stop];
            logic [RING_STOPS_WIDTH-1:0] \//@0$dest ;
            assign \//@0$dest = Stop_INPIPE_dest_a0[stop];
            logic  \//@2$empty ;
            assign \//@2$empty = Stop_INPIPE_empty_a2[stop];
            logic  \//@2$full ;
            assign \//@2$full = Stop_INPIPE_full_a2[stop];
            logic  \//@1$grow ;
            assign \//@1$grow = Stop_INPIPE_grow_a1[stop];
            logic  \//@1$out_blocked ;
            assign \//@1$out_blocked = Stop_INPIPE_out_blocked_a1[stop];
            logic  \//@0$parity ;
            assign \//@0$parity = Stop_INPIPE_parity_a0[stop];
            logic  \//@1$push ;
            assign \//@1$push = Stop_INPIPE_push_a1[stop];
            logic  \//@1$reset ;
            assign \//@1$reset = Stop_INPIPE_reset_a1[stop];
            logic  \//@1$shrink ;
            assign \//@1$shrink = Stop_INPIPE_shrink_a1[stop];
            logic  \//@0$trans_avail ;
            assign \//@0$trans_avail = Stop_INPIPE_trans_avail_a0[stop];
            logic  \//@1$trans_valid ;
            assign \//@1$trans_valid = Stop_INPIPE_trans_valid_a1[stop];
            logic  \//@1$two_valid ;
            assign \//@1$two_valid = Stop_INPIPE_two_valid_a1[stop];
            logic [$clog2((6)+1)-1:0] \//@1$valid_count ;
            assign \//@1$valid_count = Stop_INPIPE_valid_count_a1[stop];
            logic  \//@1$would_bypass ;
            assign \//@1$would_bypass = Stop_INPIPE_would_bypass_a1[stop];

            //
            // Scope: >entry[(6)-1:0]
            //
            for (entry = 0; entry <= (6)-1; entry++) begin : \>entry 
               logic  \///@1$ANY ;
               assign \///@1$ANY  = 1'b1;
               logic  \///@1$State ;
               assign \///@1$State = Stop_INPIPE_Entry_State_a1[stop][entry];
               logic [7:0] \///@1$data ;
               assign \///@1$data = Stop_INPIPE_Entry_data_a1[stop][entry];
               logic [RING_STOPS_WIDTH-1:0] \///@1$dest ;
               assign \///@1$dest = Stop_INPIPE_Entry_dest_a1[stop][entry];
               logic  \///@2$is_head ;
               assign \///@2$is_head = Stop_INPIPE_Entry_is_head_a2[stop][entry];
               logic  \///@1$is_tail ;
               assign \///@1$is_tail = Stop_INPIPE_Entry_is_tail_a1[stop][entry];
               logic  \///@2$next_entry_state ;
               assign \///@2$next_entry_state = Stop_INPIPE_Entry_next_entry_state_a2[stop][entry];
               logic  \///@1$parity ;
               assign \///@1$parity = Stop_INPIPE_Entry_parity_a1[stop][entry];
               logic  \///@2$prev_entry_state ;
               assign \///@2$prev_entry_state = Stop_INPIPE_Entry_prev_entry_state_a2[stop][entry];
               logic  \//@1$prev_entry_was_tail ;
               assign \//@1$prev_entry_was_tail = Stop_INPIPE_Entry_prev_entry_was_tail_a1[stop][entry];
               logic  \//@1$push ;
               assign \//@1$push = Stop_INPIPE_Entry_push_a1[stop][entry];
               logic  \///@2$reconstructed_is_tail ;
               assign \///@2$reconstructed_is_tail = Stop_INPIPE_Entry_reconstructed_is_tail_a2[stop][entry];
               logic  \///@2$reconstructed_valid ;
               assign \///@2$reconstructed_valid = Stop_INPIPE_Entry_reconstructed_valid_a2[stop][entry];
               logic  \///@1$valid ;
               assign \///@1$valid = Stop_INPIPE_Entry_valid_a1[stop][entry];
            end
         end

         //
         // Scope: |outpipe
         //
         if (1) begin : \|outpipe 
            logic  \//?$trans_valid@1$ANY ;
            assign \//?$trans_valid@1$ANY  = 1'b1;
            logic  \//@0$blocked ;
            assign \//@0$blocked = Stop_OUTPIPE_blocked_a0[stop];
            logic [7:0] \//?$trans_valid@1$data ;
            assign \//?$trans_valid@1$data = Stop_OUTPIPE_data_a1[stop];
            logic  \//?$trans_valid@1$parity ;
            assign \//?$trans_valid@1$parity = Stop_OUTPIPE_parity_a1[stop];
            logic  \//@0$trans_avail ;
            assign \//@0$trans_avail = Stop_OUTPIPE_trans_avail_a0[stop];
            logic  \//@0$trans_valid ;
            assign \//@0$trans_valid = Stop_OUTPIPE_trans_valid_a0[stop];
         end

         //
         // Scope: |rg
         //
         if (1) begin : \|rg 
            logic  \//?$valid@1$ANY ;
            assign \//?$valid@1$ANY  = 1'b1;
            logic [7:0] \//?$valid@1$data ;
            assign \//?$valid@1$data = Stop_RG_data_a1[stop];
            logic [RING_STOPS_WIDTH-1:0] \//@0$dest ;
            assign \//@0$dest = Stop_RG_dest_a0[stop];
            logic  \//?$valid@1$parity ;
            assign \//?$valid@1$parity = Stop_RG_parity_a1[stop];
            logic  \//@0$pass_on ;
            assign \//@0$pass_on = Stop_RG_pass_on_a0[stop];
            logic  \//@0$passed_on ;
            assign \//@0$passed_on = Stop_RG_passed_on_a0[stop];
            logic  \//@0$valid ;
            assign \//@0$valid = Stop_RG_valid_a0[stop];
         end
      end

      //
      // Scope: |reset
      //
      if (1) begin : \|reset 
         logic  \/@0$reset ;
         assign \/@0$reset = RESET_reset_a0;
      end


   end

// ---------- Generated Code Ends ----------
`line 51 "ring.m4out.tlv"
//_\TLV
   // Hierarchy
   //_>stop
   
   // Reset
   //_|reset
      //_@0
         assign RESET_reset_a0 = reset;

   // FIFOs
   for (stop = 0; stop <= RING_STOPS-1; stop++) begin : L1b_Stop //_>stop
      // Inputs
      //_|inpipe
         //_@0
            assign Stop_INPIPE_data_a0[stop][7:0] = data_in[stop];
            assign Stop_INPIPE_parity_a0[stop] = 1'b0;
            assign Stop_INPIPE_dest_a0[stop][RING_STOPS_WIDTH-1:0] = dest_in[stop];
            assign Stop_INPIPE_trans_avail_a0[stop] = !RESET_reset_a2 && valid_in[stop];
         //_@1
            assign Stop_INPIPE_trans_valid_a1[stop] = Stop_INPIPE_trans_avail_a1[stop] && ! Stop_INPIPE_blocked_a1[stop];

      // FIFOs
      `line 415 "pipeflow_tlv.m4"
         //|default
         //   @0
         /*SV_plus*/
            localparam bit [$clog2((6)+1)-1:0] full_mark = 6;
         
         // FIFO Instantiation
         
         // Hierarchy declarations
         //_|inpipe
            //_>entry
         //_|fo
            //_>entry
         
         // Hierarchy
         //_|inpipe
            //_@1
               assign Stop_INPIPE_reset_a1[stop] = RESET_reset_a1;
               assign Stop_INPIPE_out_blocked_a1[stop] = Stop_FO_blocked_a0[stop];
               assign Stop_INPIPE_blocked_a1[stop] = Stop_INPIPE_full_a2[stop] && Stop_INPIPE_out_blocked_a1[stop];
               `BOGUS_USE(Stop_INPIPE_blocked_a1[stop])   // Not required to be consumed elsewhere.
               assign Stop_INPIPE_would_bypass_a1[stop] = Stop_INPIPE_empty_a2[stop];
               assign Stop_INPIPE_bypass_a1[stop] = Stop_INPIPE_would_bypass_a1[stop] && ! Stop_INPIPE_out_blocked_a1[stop];
               assign Stop_INPIPE_push_a1[stop] = Stop_INPIPE_trans_valid_a1[stop] && ! Stop_INPIPE_bypass_a1[stop];
               assign Stop_INPIPE_grow_a1[stop]   =   Stop_INPIPE_trans_valid_a1[stop] &&   Stop_INPIPE_out_blocked_a1[stop];
               assign Stop_INPIPE_shrink_a1[stop] = ! Stop_INPIPE_empty_a2[stop] && ! Stop_INPIPE_trans_avail_a1[stop] && ! Stop_INPIPE_out_blocked_a1[stop];
               assign Stop_INPIPE_valid_count_a1[stop][$clog2((6)+1)-1:0] = Stop_INPIPE_reset_a1[stop] ? '0
                                                           : Stop_INPIPE_valid_count_a2[stop] + (
                                                                Stop_INPIPE_grow_a1[stop]   ? { {($clog2((6)+1)-1){1'b0}}, 1'b1} :
                                                                Stop_INPIPE_shrink_a1[stop] ? '1
                                                                        : '0
                                                             );
               // At least 2 valid entries.
               //$two_valid = | $ValidCount[m4_counter_width-1:1];
               // but logic depth minimized by taking advantage of prev count >= 4.
               assign Stop_INPIPE_two_valid_a1[stop] = | Stop_INPIPE_valid_count_a2[stop][$clog2((6)+1)-1:2] || | Stop_INPIPE_valid_count_a1[stop][2:1];
               // These are an optimization of the commented block below to operate on vectors, rather than bits.
               // TODO: Keep optimizing...
               assign {Stop_INPIPE_Entry_prev_entry_was_tail_a1[stop]} = {Stop_INPIPE_Entry_reconstructed_is_tail_a2[stop][4:0], Stop_INPIPE_Entry_reconstructed_is_tail_a2[stop][5]} /* circular << */;
               assign {Stop_INPIPE_Entry_push_a1[stop]} = {6{Stop_INPIPE_push_a1[stop]}} & Stop_INPIPE_Entry_prev_entry_was_tail_a1[stop];
               for (entry = 0; entry <= (6)-1; entry++) begin : L2b_INPIPE_Entry //_>entry
                  // Replaced with optimized versions above:
                  // $prev_entry_was_tail = >entry[(entry+(m4_depth)-1)%(m4_depth)]$reconstructed_is_tail#+1;
                  // $push = |m4_in_pipe$push && $prev_entry_was_tail;
                  assign Stop_INPIPE_Entry_valid_a1[stop][entry] = (Stop_INPIPE_Entry_reconstructed_valid_a2[stop][entry] && ! Stop_FO_Entry_pop_a0[stop][entry]) || Stop_INPIPE_Entry_push_a1[stop][entry];
                  assign Stop_INPIPE_Entry_is_tail_a1[stop][entry] = Stop_INPIPE_trans_valid_a1[stop] ? Stop_INPIPE_Entry_prev_entry_was_tail_a1[stop][entry]  // shift tail
                                                     : Stop_INPIPE_Entry_reconstructed_is_tail_a2[stop][entry];  // retain tail
                  assign Stop_INPIPE_Entry_State_a1[stop][entry] = Stop_INPIPE_reset_a1[stop] ? 1'b0
                                             : Stop_INPIPE_Entry_valid_a1[stop][entry] && ! (Stop_INPIPE_two_valid_a1[stop] && Stop_INPIPE_Entry_is_tail_a1[stop][entry]); end
            //_@2
               assign Stop_INPIPE_empty_a2[stop] = ! Stop_INPIPE_two_valid_a2[stop] && ! Stop_INPIPE_valid_count_a2[stop][0];
               assign Stop_INPIPE_full_a2[stop] = (Stop_INPIPE_valid_count_a2[stop] == full_mark);  // Could optimize for power-of-two depth.
            for (entry = 0; entry <= (6)-1; entry++) begin : L2c_INPIPE_Entry //_>entry
               //_@2
                  assign Stop_INPIPE_Entry_prev_entry_state_a2[stop][entry] = Stop_INPIPE_Entry_State_a2[stop][(entry+(6)-1)%(6)];
                  assign Stop_INPIPE_Entry_next_entry_state_a2[stop][entry] = Stop_INPIPE_Entry_State_a2[stop][(entry+1)%(6)];
                  assign Stop_INPIPE_Entry_reconstructed_is_tail_a2[stop][entry] = (  Stop_INPIPE_two_valid_a2[stop] && (!Stop_INPIPE_Entry_State_a2[stop][entry] && Stop_INPIPE_Entry_prev_entry_state_a2[stop][entry])) ||
                                           (! Stop_INPIPE_two_valid_a2[stop] && (!Stop_INPIPE_Entry_next_entry_state_a2[stop][entry] && Stop_INPIPE_Entry_State_a2[stop][entry])) ||
                                           (Stop_INPIPE_empty_a2[stop] && (entry == 0));  // need a tail when empty for push
                  assign Stop_INPIPE_Entry_is_head_a2[stop][entry] = Stop_INPIPE_Entry_State_a2[stop][entry] && ! Stop_INPIPE_Entry_prev_entry_state_a2[stop][entry];
                  assign Stop_INPIPE_Entry_reconstructed_valid_a2[stop][entry] = Stop_INPIPE_Entry_State_a2[stop][entry] || (Stop_INPIPE_two_valid_a2[stop] && Stop_INPIPE_Entry_prev_entry_state_a2[stop][entry]); end
         // Write data
         //_|inpipe
            //_@1
               for (entry = 0; entry <= (6)-1; entry++) begin : L2d_INPIPE_Entry //_>entry
                  //?$push
                  //   $aNY = |m4_in_pipe['']m4_trans_hier$ANY;
                  assign {Stop_INPIPE_Entry_data_a1[stop][entry][7:0], Stop_INPIPE_Entry_dest_a1[stop][entry][RING_STOPS_WIDTH-1:0], Stop_INPIPE_Entry_parity_a1[stop][entry]} = Stop_INPIPE_Entry_push_a1[stop][entry] ? {Stop_INPIPE_data_a1[stop], Stop_INPIPE_dest_a1[stop], Stop_INPIPE_parity_a1[stop]} : {Stop_INPIPE_Entry_data_a2[stop][entry], Stop_INPIPE_Entry_dest_a2[stop][entry], Stop_INPIPE_Entry_parity_a2[stop][entry]} /* RETAIN */; end
         // Read data
         //_|fo
            //_@0
               //$pop  = ! >m4_top|m4_in_pipe$empty#m4_align(m4_in_at + 1, m4_out_at) && ! $blocked;
               for (entry = 0; entry <= (6)-1; entry++) begin : L2b_FO_Entry //_>entry
                  assign Stop_FO_Entry_is_head_a0[stop][entry] = Stop_INPIPE_Entry_is_head_a2[stop][entry];
                  assign Stop_FO_Entry_pop_a0[stop][entry]  = Stop_FO_Entry_is_head_a0[stop][entry] && ! Stop_FO_blocked_a0[stop];
                  //_>read_masked
                     assign {Stop_FO_Entry_ReadMasked_data_a0[stop][entry][7:0], Stop_FO_Entry_ReadMasked_dest_a0[stop][entry][RING_STOPS_WIDTH-1:0], Stop_FO_Entry_ReadMasked_parity_a0[stop][entry]} = Stop_FO_Entry_is_head_a0[stop][entry] ? {Stop_INPIPE_Entry_data_a2[stop][entry], Stop_INPIPE_Entry_dest_a2[stop][entry], Stop_INPIPE_Entry_parity_a2[stop][entry]} /* $aNY */ : '0;
                  //_>accum
                     assign {Stop_FO_Entry_Accum_data_a0[stop][entry][7:0], Stop_FO_Entry_Accum_dest_a0[stop][entry][RING_STOPS_WIDTH-1:0], Stop_FO_Entry_Accum_parity_a0[stop][entry]} = ((entry == 0) ? '0 : {Stop_FO_Entry_Accum_data_a0[stop][(entry+(6)-1)%(6)], Stop_FO_Entry_Accum_dest_a0[stop][(entry+(6)-1)%(6)], Stop_FO_Entry_Accum_parity_a0[stop][(entry+(6)-1)%(6)]}) |
                                {Stop_FO_Entry_ReadMasked_data_a0[stop][entry], Stop_FO_Entry_ReadMasked_dest_a0[stop][entry], Stop_FO_Entry_ReadMasked_parity_a0[stop][entry]}; end
               //_>head
                  assign Stop_FO_Head_trans_avail_a0[stop] = Stop_FO_trans_avail_a0[stop];
                  //_?$trans_avail
                     assign {w_Stop_FO_Head_data_a0[stop][7:0], w_Stop_FO_Head_dest_a0[stop][RING_STOPS_WIDTH-1:0], w_Stop_FO_Head_parity_a0[stop]} = {Stop_FO_Entry_Accum_data_a0[stop][(6)-1], Stop_FO_Entry_Accum_dest_a0[stop][(6)-1], Stop_FO_Entry_Accum_parity_a0[stop][(6)-1]};
         
         // Bypass
         //_|fo
            //_@0
               // Available output.  Sometimes it's necessary to know what would be coming to determined
               // if it's blocked.  This can be used externally in that case.
               //_>fifo_head
                  assign Stop_FO_FifoHead_trans_avail_a0[stop] = Stop_FO_trans_avail_a0[stop];
                  //_?$trans_avail
                     
                     assign {w_Stop_FO_FifoHead_data_a0[stop][7:0], w_Stop_FO_FifoHead_dest_a0[stop][RING_STOPS_WIDTH-1:0], w_Stop_FO_FifoHead_parity_a0[stop]} = Stop_INPIPE_would_bypass_a1[stop]
                                  ? {Stop_INPIPE_data_a1[stop], Stop_INPIPE_dest_a1[stop], Stop_INPIPE_parity_a1[stop]}
                                  : {Stop_FO_Head_data_a0[stop], Stop_FO_Head_dest_a0[stop], Stop_FO_Head_parity_a0[stop]};
               assign Stop_FO_trans_avail_a0[stop] = ! Stop_INPIPE_would_bypass_a1[stop] || Stop_INPIPE_trans_avail_a1[stop];
               assign Stop_FO_trans_valid_a0[stop] = Stop_FO_trans_avail_a0[stop] && ! Stop_FO_blocked_a0[stop];
               //_?$trans_valid
                  assign {w_Stop_FO_data_a0[stop][7:0], w_Stop_FO_dest_a0[stop][RING_STOPS_WIDTH-1:0], w_Stop_FO_parity_a0[stop]} = {Stop_FO_FifoHead_data_a0[stop], Stop_FO_FifoHead_dest_a0[stop], Stop_FO_FifoHead_parity_a0[stop]};
                               
                               
                               
         /* Alternate code for pointer indexing.  Replaces $ANY expression above.
         
         // Hierarchy
         |inpipe
            >entry2[(6)-1:0]
         
         // Head/Tail ptrs.
         |inpipe
            @1
               $NextWrPtr[\$clog2(6)-1:0] =
                   $reset       ? '0 :
                   $trans_valid ? ($NextWrPtr#+1 == (6 - 1))
                                    ? '0
                                    : $NextWrPtr#+1 + {{(\$clog2(6)-1){1'b0}}, 1'b1} :
                                  $RETAIN;
         |fo
            @0
               $NextRdPtr[\$clog2(6)-1:0] =
                   >stop|inpipe$reset#+1
                                ? '0 :
                   $trans_valid ? ($NextRdPtr#+1 == (6 - 1))
                                    ? '0
                                    : $NextRdPtr#+1 + {{(\$clog2(6)-1){1'b0}}, 1'b1} :
                                  $RETAIN;
         // Write FIFO
         |inpipe
            @1
               $dummy = '0;
               ?$trans_valid
                  // This doesn't work because SV complains for FIFOs in replicated context that
                  // there are multiple procedures that assign the signals.
                  // Array writes can be done in an SV module.
                  // The only long-term resolutions are support for module generation and use
                  // signals declared within for loops with cross-hierarchy references in SV.
                  // TODO: To make a simulation-efficient FIFO, use DesignWare.
                  {>entry2[$NextWrPtr#+1]$$ANY} = $ANY;
         // Read FIFO
         |fo
            @0
               >read2
                  $trans_valid = |fo$trans_valid;
                  ?$trans_valid
                     $ANY = >stop|inpipe>entry2[|fo$NextRdPtr#+1]$ANY#+1;
                  `BOGUS_USE($dummy)
               ?$trans_valid
                  $ANY = >read2$ANY;
         */
      //_\end_source
      `line 72 "ring.m4out.tlv"

      // Outputs
      //_|inpipe
         //_@1
            assign accepted[stop] = Stop_INPIPE_trans_valid_a1[stop];
      //_|outpipe
         //_@2
            assign data_out[stop] = Stop_OUTPIPE_data_a2[stop];
            `BOGUS_USE(Stop_OUTPIPE_parity_a2[stop])
            assign valid_out[stop] = Stop_OUTPIPE_trans_valid_a2[stop]; end

   // Instantiate the ring.
   `line 643 "pipeflow_tlv.m4"
      
      // Logic
      for (stop = 0; stop <= RING_STOPS-1; stop++) begin : L1c_Stop //_>stop
         //|default
         //   @0
         /*SV_plus*/
            int prev_hop = (stop + RING_STOPS - 1) % RING_STOPS;
         //_|fo
            //_@0
               assign Stop_FO_blocked_a0[stop] = Stop_RG_passed_on_a0[stop];
         //_|rg
            //_@0
               assign Stop_RG_passed_on_a0[stop] = Stop_RG_pass_on_a1[prev_hop];
               assign Stop_RG_valid_a0[stop] = ! RESET_reset_a1 &&
                        (Stop_RG_passed_on_a0[stop] || Stop_FO_trans_avail_a0[stop]);
               assign Stop_RG_pass_on_a0[stop] = Stop_RG_valid_a0[stop] && ! Stop_OUTPIPE_trans_valid_a0[stop];
               assign Stop_RG_dest_a0[stop][RING_STOPS_WIDTH-1:0] =
                  Stop_RG_passed_on_a0[stop]
                     ? Stop_RG_dest_a1[prev_hop]
                     : Stop_FO_dest_a0[stop];
            //_@1
               //_?$valid
                  assign {w_Stop_RG_data_a1[stop][7:0], w_Stop_RG_parity_a1[stop]} =
                     Stop_RG_passed_on_a1[stop]
                        ? {Stop_RG_data_a2[prev_hop], Stop_RG_parity_a2[prev_hop]}
                        : {Stop_FO_data_a1[stop], Stop_FO_parity_a1[stop]};
         //_|outpipe
            // Ring out
            //_@0
               assign Stop_OUTPIPE_trans_avail_a0[stop] = Stop_RG_valid_a0[stop] && (Stop_RG_dest_a0[stop] == stop);
               assign Stop_OUTPIPE_blocked_a0[stop] = 1'b0;
               assign Stop_OUTPIPE_trans_valid_a0[stop] = Stop_OUTPIPE_trans_avail_a0[stop] && ! Stop_OUTPIPE_blocked_a0[stop];
            //_?$trans_valid
               //_@1
                  assign {w_Stop_OUTPIPE_data_a1[stop][7:0], w_Stop_OUTPIPE_parity_a1[stop]} = {Stop_RG_data_a1[stop], Stop_RG_parity_a1[stop]}; end
   //_\end_source
   `line 85 "ring.m4out.tlv"

//_\SV

endmodule


// Undefine macros defined by SandPiper.
`undef BOGUS_USE
`undef WHEN
